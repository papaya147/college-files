module testbench;
  reg [0:15]x;
  reg [0:3]s;
  wire f;
  mux16to1 sto1(x, s, f);
  initial begin
    x[0] = 1; x[1] = 1; x[2] = 1; x[3] = 1; x[4] = 1; x[5] = 0; x[6] = 0; x[7] = 0; x[8] = 0; x[9] = 0; x[10] = 0; x[11] = 1; x[12] = 0; x[13] = 1; x[14] = 0; x[15] = 0;
    s[0] = 0; s[1] = 0; s[2] = 0; s[3] = 0;
    #100
    s[0] = 0; s[1] = 0; s[2] = 0; s[3] = 1;
    #100
    s[0] = 0; s[1] = 0; s[2] = 1; s[3] = 0;
    #100
    s[0] = 0; s[1] = 0; s[2] = 1; s[3] = 1;
    #100
    s[0] = 0; s[1] = 1; s[2] = 0; s[3] = 0;
    #100
    s[0] = 0; s[1] = 1; s[2] = 0; s[3] = 1;
    #100
    s[0] = 0; s[1] = 1; s[2] = 1; s[3] = 0;
    #100
    s[0] = 0; s[1] = 1; s[2] = 1; s[3] = 1;
    #100
    s[0] = 1; s[1] = 0; s[2] = 0; s[3] = 0;
    #100
    s[0] = 1; s[1] = 0; s[2] = 0; s[3] = 1;
    #100
    s[0] = 1; s[1] = 0; s[2] = 1; s[3] = 0;
    #100
    s[0] = 1; s[1] = 0; s[2] = 1; s[3] = 1;
    #100
    s[0] = 1; s[1] = 1; s[2] = 0; s[3] = 0;
    #100
    s[0] = 1; s[1] = 1; s[2] = 0; s[3] = 1;
    #100
    s[0] = 1; s[1] = 1; s[2] = 1; s[3] = 0;
    #100
    s[0] = 1; s[1] = 1; s[2] = 1; s[3] = 1;
    #100
    s[0] = 0;
  end

initial
  begin
    $dumpfile("dump.vcd");
    $dumpvars(1);
  end 
endmodule